DBCDL40 COPYRIGHT � 1997-2002 DATA BECKER GmbH & Co. KG       հ   �   �  �  s  #  s  �"  s  	&  S  \)  S  �,  �T  `�  s  Ӈ  s  F�  s  ��  �  l�  �  �  �  ���� JFIF      �� C 


�� C		��  � �" ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ���x�`�i�Ha�K��0UU$�z ;ׂ�\��Ǉ��A��Ζ�j�X�VF`fxٻ	��	q���F��@��b��c�Q���׼W������R9��KX�i���
:T����W�k� ����h�J*O�1%��-��}ǁӞ>AOx��?���i��$�����XI�i������hv�}z�{�|�=_�|�/5�7jmEyj�f��>6���$�^����c#�iM�q7U�I��$� ������!�x�J��__xfW�"y.u9�)�'XYv�e���J�;y����������2\�"u
Y��A
A ��j��4�=~��k�[]��|����H�%�B�+����|tԕQ����N*.J2�ݷv�h?�N��x^�R/6���WL���j����;�E��U� �����L�^���������K������d9`$dd�p�@<�[~�zV�6��6��Dig�Ӯ��[�pѳ2ªdR��=��p^$�k�x�����-�[^[	␆Qr���9���,�08�k'�i��ǝJ^��O��3�XEy��X^æ_�(�2�	��qZ2�I�� ��ǯ�G�w��i�;�*�� ˕���]Hn���g��k�j:��{8��Imⷁ�Egfy�W�LF
'�Y7 �Yv� �G�?Bu���,&u���3���]H9!s6J��k2	9���^ܬ롙�!+_�y��?J�����{�������� L`�s4C )$}����98�����S�K�;���;&�ã`��� �¼J�z�wi����q��q�7�n��QEr��Q�<V�I4�$0ƥ�I*���I= �J��?��#��?o,�Dʫvm��I�g������s�Npgz]y�#�����/��8�W�����mtKW�EY�$vb�']�M�",�F�w�\/�[xoU�5o�9��N��0�麊�A#�*��>�Kn�.�j�A�� ��{MrV��+I=�����th�a'G���(�id,U]�}e*1�yc��5�3�>yk'�Yv����1I�*�(,ŏ��O��QEuc������D�4.�:������V��6����OZŪ�ơ3i���KǺ'����%���Q��O�)� �|ua}u"�mm���� ��HI$� �q�z�>-ҵby�n�n>�!�[S<�Q#B�2JĀ�.P���FG�f�Ɗ��Y�OA�V�K�+7�&�ǧ|+�ym�j�}?E�Gڻ� ��<O��w|fdo0 [��Ӄ����1�`��O
�O<v�t�����9. �J�q�ZY̮XG��N��
䫧)�/����:��ɻ��j��VV��m'_�$Ԭ!�t]���)�ˏF�ã dZ�W�4���&֨�a��~�W70"+p������(~�21;7��凩|��{�Aܐ��EԎ'��_1kB�.rp�?�a�W	�I�f��[�ۖ͝����*�/�)��a`*�ʠ�,]�o�$��L�VP��=$��=+U��4�/�'K�I�|r�B?� �� �V��_���ܹ�t���V
��?/m#��rf ܝ��;�����Pt'�ӡ��<Tqt���F��Ǟ+�����ܡ�e�o��JxQ����@9�����yh��)#���7W&!���g͍��+�!�p�?H~����6��(����]�L�����~R#�{|����ڇ��uGX����[��n�q�*A#���
��\J*��/�����-$���#�s\G=g/�o_�C����4{�-�,�جŶ�I�'�� � j��A�\��T�����\�񰺄e�+�0� W��Ҳ��Jg�(�:;�=�|nc]��Fx�����۶�<����5���mn�O����3�� �.#�X�F&F;Hݿ m?(���ѼAb����&X��'ߦ�D��3�`�`8㞃��oȮD����GU{jom^���-��2�k+��?,кH��v��$�ERӴ9��B��/x�i-�I�+�j�09RY"��D8�YXdA"��o�G,���;�ax�Y5H٤fVh�����P�˒I<C&�4o��(�O��ƸIs� 
NI���X�S�����tӕjk��F��2;�+I�ѵk=F��^4���d��n�a��DYX0�,�.@�:�a�A�ѯ<��횺yb�+�f����_2T�H��Ky����$ Y�W7O�"�4F��in���+� Rd��8rS�#oK
��V��m۽��zU�hv��,����H�r�>�(�v3�T}�ˎ[$��-���Iip]�is4~Tq�k(�6��	�$��A<��ּϷ�s�%��?�;*���.���ԩ#���ɷ��M���I�9E��߲��{� �x ���h֗�ZzC}��tٮ|��p.J����H_}�<�i��%��N� y�x-oF�&��\X�t�dy�VW��W3�!�䫀�K�(ȯ�>x�q�t��DmRռ���.��_h<���𷌼5yw�-W���n�]�do*�I-(��;�7d]�YFpH?C���&{oLz��-Ȓ12�� �y� s�����(�їx�S�˱�":�=�C�k\��j��u-����O�e�[��FHʢ�e$)�n�F��9����S����ޭu���4�=�,eU�64X�͌� �i~Қ���x�d�M��s�\^Z�jZ8�%d��$�1�덠��F;+{x� �cX��B$h0��` ; +��me�$y���''�m��QE�pGqm�-�$�62�(e89qRQ@��0ga���p�&[��*;�h7n^}N���i-#bx#��$~&���� �� ���7wv)s�αܼ������T�ORFO`8�5ᇍ�s���j�&�d�g��xkG�X%�J��H3�۠1川�e�n;�֛'��Ya��`���kd+��c��Wٞ4�m�x���'���P���Q9X)c՗'�� ���[Y�h��b��U�����8lD1)�Y���:�).i]=�N�N�ӖE����es#�c� ��S�9�b�+���
(��9�xsA�#�U׭c��ҡ�V�h���eA}����� ���n|1�Ւ�Xk,sGo�\ �mj�B���@*7ѺTZƜu}6{?��j&ZH�7;r7.���S�<���6�M�%[�Ԣ�w�� ]��'>J"��$d�k7�[Fo���lb|v�
����siw�YOtQnlD���.�n�71���[8��;H�bgY&
�)Uf�$N{d�M[��/�7�^�>� ��^�6�H�(�^2���v��������n�O��@�#����;���ܯ=�~������b�q����K4QEnrU}B�*�{˗1���I)m�I��@nX��>x��ƾ��.|�B�;�e
�.9m���A �;pA����2kO,��Gړ�lmz�ˁ������=3P�z���]E/�``_8�dn� �p�C��G�����M���>��?��� h�jZ��T	ª��7dQݎ?�8 �����}N�����˛�Y_ nf9'���Y�<��5K�s����@�n#2��26(����{� Uy|e�@��֟��)�Q�B��
�#�3�N2~��/��6KݲF�����n'����̢H\:��U�G}"��@�(���O�xoT���)���H�)�)&T���g�Cg9�k�6�{�h��W�Ku,�hk��M��Ѡbc=0F��ۜ�I7>%����:�ΐ_Ou0ﵖ�1-ФH�p��Y��G��+���Q�ѽ֥�,r��HF��w`c9��+&��w��J^��f�q���ISU�uq���h�C�X��z�v�� `���w�<a�j�/6���V���kW��+E�"W̍��0���2uO�/��� ���v1���� �-y� ��P>`Yrx�ھ
��sy��F���."���c�u�#�.CJ�o
5R	��$y�*��R����e�pķm'��_�;�*;k��-�C*GH�?�V�u4�=�b�����|�q�`��=�'��:ױ}.|�voT�Cѯ�)Q����K�D��K=��6?�'�.�ۓymx��	k�|��U	�6�~q�N��䜍��߇�ܭ����#���$��\��N�o�#x���jXx�mB���G�kCrΊ�PXʫ6�$*���%���7�� �0�^�o��z��O y�����z��r\y�1Y"#�0\L�$�'����)�lK��a�n�v��u�K��!�kXw;�2F�b1��e�\��|������r�o�.<'�E:���C�8�NA g���\>8b$)��vB���s�#s����׮x�_��Wm�_�q����?x���M�Z[�\�<�_�NB>a�E��n�[0����v�#؋���*As��DN|����� ���t<Z�V�d��V��zRI�m�1_$I��r\3�����x"�j�n4ԅ��Ϙ�J�l�Twc�<�|�� ����������<��5�g�O�K��V����cc}�������#�%�pH�Mv��m����a�,`��sF�4�k N�S�#*A9�^=xm�/보Oyb�Č��睁r݆�瓅��ݬ���:��ʈ� �4�YU�pHQ��99S�z�6��OC)EIi?S���-7ǳ_܈��:岴�$��P���#��$�qZ�/�$�</��C�y�ۻFbM쯌)��8$��'�kNd��9$��9?��	-��M�r���1,@'�6}�D����3��uʓ��~����<n|o�(`���ݱ_����X�8^������τ�7��v�,��[Z�y#Y���A<%���2�?!
��:���/��/�������Yc�Ѡȍ���@~|�����:���e�\Tb�k�_���g���1��:+�:Iiƭ�[���.ߗ<��ų��?I��0jv7w)�[\F�J�#r���j��=wB|�:�]��,U'��?3�g@�W�F�a�ޱ�V�q�on���f%�vnQ呈�5)�nkҫ����n�y2̶Wq���<K'w��c�ldT���g�[�!���.}NKx��{�h�g�j��|���!'���ݘ�j��u"�x��kQ������~��QU4�V�Z�[���$OPpAA�5n�w8ڶ�(��QE Q\��|u��Ea��k���)�FJ+8�V`�&nf,0��&�U�Q���:Y�X"y1U!�� �?A^w���S�H�෵���m�g�K�& ���yxb
����pz�e�k�5����PG�ľ}�ݓ�X��Ml����ub�libp�;����k�ߍ>�R(�y׷�X�f��.xgm�(<�ğ�Մ��\��Q�
mIF��cC�q�]�k?هY� L��\��Õa3,��	7��#$���U������%��bZ�)U�sI$��I'�9��iW��k��E���,"�ӳ������QE�zMWJ��4��/�K�I�d�?B?�� _5�^�����.��k:d�I�]�V�&Ƥ|�O�?/?t1�~�ꡈ���ۡÊ���G���ks��[YxJML�"�w�<xnAmΌT`y��N8V8
���g���ig�;)����
���$�j�`�t����F�_
�u���6�㇒�T{-Q�yV�!w��#Ѱ�n�o�� �V�ow͜v:��y,sŕ���}8rO���c(Զ���c��帊-��������ߊ��]�wr=�Zζ�\9M�V��	�1�g9۴���㏍��2�����j������=���Ϛ�!��r���c�WU�O������t[���m�:��NUU�9��!a��1ǃ��u��m�.t�[�,v����+2
��ێs۶+��n-ye�A�4��s��I���ڥ�7��>�%�,�����-�w�U��)�������%�^��bw*d�ln�Ԏ�Vn��E�5��k�����;�,n��-Ք���"���0�ii���vYm��Zb�\�B��%��!1���U炲9��75}�B�7d�ف�x��:����[,$�qiu;ۙԌ����$So���a����/<C��|L�u+Y���[��)]����fFtm�~Wl�=�@��|Iyu)���F��F�I$Wy8
X�P>b;�zǂ~	h�����mJ&��6�pV0O8#�-ʂ1\5q�i��s>����P˱5��9Ww���3�������|mf�?�!�Q$*��Wjħ�
����g�?Lh�|-�.�--Cؤ�X�$�I=I� �iQ^#<C�E���&�^:��aEW������� JFIF      �� C 


�� C		��  � �" ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��(������ JFIF      �� C 


�� C		��  � �" ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��(������ JFIF      �� C 


�� C		��  � �" ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��(������ JFIF      �� C 


�� C		��  d �" ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��(������ JFIF      �� C 


�� C		��  d �" ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��(������ JFIF      �� C 


�� C		��   " ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ��( ��( ��( ��|C�'��V���6���]� �Q�ln�8�5�/��oo7A��_������U�?t�� �vA�]Tp�k�N�N6�~�Z�[� ^���_�i��syq��c|ӸD\��������w�?����dseU8��T0<�#��~r��I�x�7S�./�3:��%P��ڽp8 �f׳K,�֣����ʒv�/=_���ǩ�Қ��W�v�ik���j����۳�s����q���"j�3GkT�Rp:rI����#����?����Twu�O��� ��Ŀ�0��/� Tu={S����F�� �ϗ���M��q��g�F��B)�#�Ԝ���oMկ�i�m>���f]�KiZ6+�q�G�j�� ��Ŀ�0��/� Xu�W��#���W��i�]*�]KƱ��7�./�]Iqg�]�2<�Hw[��A�NV<�����[:����oB5*{��m���}��[AI��H� 2A� c�(I>���W���z�S��4�+�v�%�<,#���c<c�.�M�/��ZѼ.�V���;-�umf����H��b�爪$R�i�g
��f�ֿ��?��� ��v�_�"�?c�/�2�H�L3$�)%�����_3c�0��J���T18�v���K�}���v��A�gPڷ�w���v�/2=�eT�X�8%G�J�=7V��`i���{�U�-�Y6�A<��=��O|G��{w�O�"X�E��^HD�����c��\� ��]v��_hӴ�}�Ō̻�ҴlW � �2��<����Jߊ=Y�jO��o�3�+�_
~кƝ8�\�5kVl�cU�h�#� V 8 O���<�<g }2�$�.絓�>r����2��My��hk%�t}C����AEW�Q@Q@Q@Q@Q@Ug\��=bך��VV˟�V��v��̀pI��M�!6��ݑjyⵂI��!�5.�H�UT�I� �^1���6�_>S����
�cS�XՆތG�#����2���$ܰ�����S�Fv�?�@5�~0��.-K_���Ӥ����<N���6�2��!l1ʠ$�"����=����fm:��X_�����O?�}'[�u�{�~+�_L�����|K��gV/����FC�e���|O����b����ޢ�g����iqq�;���n8���?<Y��x�F�>"jwR���X��Þ(�f�l+R�4�A�v�Y.,�g�VQ#�	1�r�S��ᆻ�_�,�[x�ƚu߈���#\}F���Ù��n��!� C���<�9�Y��7��\����� ���~�kJZ�����ӻ>���+���+�?g�Mֿ�� �4�[� +��>�
ɳ>fq�g�kUTi��^�V���T��� ���^��������i�i��uW�tr�x�9b0A��<N8���c���zm��&vZ��4���#m�EP��l0ۺ y<�!���p�z����L��y/,n ��[e��.�d����YK�r���#���֓�v�sJ����麶����]_Iiq��R!ڨ�c�y؀|�ꟈ慢X6���:T%Ė1ʷҳ���@
��0�<c�]|�=5/��3G��-��,�[�R�����T�9-zz*�|����3�/x�Z�|.�V����.ot�f�����8��e�h���<Q h�xd��e�1�ǅ�G�[O	O���u/�/�m���
�+A�Q��bd�m�i_pl6VY")���J�������X�!�pi�[]z����������2���� �_c����g��T�fL�S<p��I�.���y�3��	$� ���k�Y�b�ľ����O_�|]n���k
IxL�*gfh����P�����	|94:R���j]"9��d�'k�:I&"���R���%GF+�)��x�Ŏ��� l�����ȼծ緆+�Wj�V����E�B��F|�y7�/�{9ů���tt�jrR�߆�m��o����/��Oğ
�~ Xe�t�*�x�R��r[�$�]��J�%��K��Ǩ��A<���42<3F��Hث+�A=����:��~��-CJ��:E��x��wL��jZ����[�^K	�}��Mlȃ>cC��i\���J� ��
����K_[C���;�"X��,Zr����"�&�N�s��P�+%5����&�r�-����<�>��}��[�O�({�tU�;�Դ��fQ��`���|��׸�Z����Aa:\�N��:�9A�K�~$��tm~�%��U����"��C H��#=�z�~&j� �E�	ua3��bv���R>�`c<��X�j.z:?���y��e��w���֊�𿋴���w�]$��i!$y���s��q�H�k�e�%f}�e�J.�QRPQE QE QEQ�5�oh����l����� �E n' �H�m�	���>:�֟�=�^6w���+a�oOen��~c�׎�k���P&V��[)
�{���w�  x��Z��5�yx|�+oh���}=��e��  ��z?ƿj��7�|?w�Kl�%����wnF� �Xɕ!�8F�"����dmo��a���4���h����g�������չ��ύo��_��Ɖ}g,w2�k�#�Y�� �aс+����2�vW�|9������4�T��F��kk'�`�6��ڪ��Ep�vm���w C,�?Ý�ƺ��K[�΅<o���nt�[=Bl��ಞ&W�a�Of�`o-��|��(��D�,�9�ç����n gffb���K;�fv%����$��u}��|���┣����_���8�;�k������y�"Ӷ��g�.5�9پ�%�TGi�Hc�Ta�8�,�Z(��G�YU&�K��QVf���,t\Xkȡ���@����>�����h�����Z��� ������ʿ�!�����h��mu?G��^\N�󰔳#:���ͩ��9�q��~�V�]�|S��l^�71l�֥[� ���*��}�p�#$�^�m���K�ɼ��,�خ݌��o�J��L�AHS���ງ��|A���ψ�ޡ�TI���#;-�� �Ŏy 9
>S�G�Ɩ�?[�Z�;Q�_�KV�}l���~C�;|>�-5����]y��77�\6#��*�"vo�!����c����mc�>6_���uj*VY�$��s�;Y%\����9~^�	�O�(�����<�mi|�E"~�"N��[W�|�����E����.�u�����G)��BD�����Uˢ��Yb����-�}� ��>i��+��0��(Ş	�|qoe�e�ı��e��m�7�eFF]VG*��[k)�G��k�N��k���$���a�갇�Ғ�ص���
�V����&�0������Vr�;�F��S���,���r�+��-�"�X@��\K#�qEY�GDQ���2F�~%��בhz����b�]�-����w�nE�ܐa�h�Kyo��U�]ۿ	���~���o�[I���Y��W8k�6o�n�6�y {��� �~�txb�J��w�4?�^��R���{}:xf�{������7����><�!�)�q�ii�^_���Ӝo_���n�ۯ�>�>��bKM�ʝ8enRE�;���#_N|;����A��F�b�aɖ��q۞N�������-�:׉tǸ������o��Qe���"�[���7�)cLD�K��D{�k��1�}C��:��7�:p�ܤ��wS��F��xb���u;0x��	���{���u��[x�öڭ��^fVX�h�pT��� ���ݯ��\��G�Bq�8��QEIaEPs��M4�1�w�F
��d�O@z����ď�Nu���IF�k�H�	��˷ y�]��㤊�|/jwK.ɮ�2��V29!�
ݰ�q�'��qm��ï�_�j�d(��N�L�p��q"nbN��3���H�B>ާ�ӹ��2U'�Z_?7���P�������h~9�-�V$h㵊���h����ne�:��~_#�Xֵ?���~� �h��t~#��y��8��K�T\$����� ���r�^������=#I�D�<i��B;]WD�F�|��#N��pG֒;��8[aty�rTB� @&�a�ͣ�7�$Qj֑��5�1Iu`e@$E�Kb>V��u#�+�i�6�������K[���Ko}�ƭQ]��QE QE ��o��_��� �k�+�>x�|!��k\gk�-a3J[��#q�d}GZ��� �K�����"玧����#\�ݎ��ǒZ�5�ƹk>���Jײ��$Q�\#Z_�_5z�k���-;J�u1���Yk�S|6�0�i�\�ԕpX7�[`?�8�87�O\xsU���ž!���F1xL�H����F��n{��r@�$h�(�_��K�3�-5��	%��>X�Nb �����g���|R�Տ��3�ί
�7N<��mn�O�����_�>+еF��Ǎ��"k��M|�6ؙgu��c�P9������R���:΀�΍��Z��DIV(̌�����'����8�Q^5���߅P�^�ڕ���[�go�i?kxc�^S��q"���`+C�O��l~#i�]޿�kIv$�?i��ءi�<���lfa�&�s�RѤar�akVkY;�ޑ�}�q�QE~�~QE QE ����ƙ��*�[��}��]M�+���pc+�t����,�p U�RVeFN�;�qᏃ�F���Z׍<A���7��TxUm�@����Cs6�8	$'3n˷W�x�E�u��'M��к�޷2Z����"0W��U1,�H�%��%q�O����>�t�-F]���kX53�Z��U�p�w)!�9GZ��x�¶~���#?�t-jK?�^�7�����e#��c�EfXI,����A��~yIQ�-?���G\ �	��^�����mc�7����wy�M>_���6�^ppxܤ�t�2��J�m5�:�	���u��Џ�A� � ����ŷ��o��P�o4��4��;T�G=���v�#+#���̬�)�� ��I��x~���P�}���V9����N�z� ���?�Ua��W��������]��O����z(��l�@��x�
xv� V�㶌�L���
� �,@�8�kZ���|_��R�ð7��qs�YY~A��9��Z��Q��T:u�8q����*�v^�֧���O��\^\��sq#K+���$�p9=��<[���x��_x�U��Kqy��j�J��7+�;KYJ�!��Y�]�I��~��=/�J�ѵi���&�:�y�����<�4J���P�C(�?�]�=#Y���o���kZ%��s�,u��E�L��T̆�6u��\#DT�E���S�T�?��3�S������Wϵ�w{��᥿��=f��c_�n5mLCu4��y�y6ƮB������A�(8��Eo��#�ss���
(�����( ��( ����k��3����}�j���'�ݷ;<�*�������q�4訩N5b�5tͩU�	��ݚ6?�w|j� ���� �$o�iN���5=O�Rb)l��Đ�G<R,�/��j8�
|̌X�(��W�0�����=�\g�������[u�~���o�iV���m�k)u=S��zts�\��xf�	��0ީ+j.��(�	V�9EP�� /�� �?�q���/�
(���$(�� (�� (�� +ʼQ��C�^��|E�K�/;M���qo$M]7��x`�^>0�nҪE�GU�t�w��Zu���;����T/�:gd����8a�����y��iϑ��������uO�-r�Tסx�T���c{v�G�ma�9d��2����|���+^9�xS���_�-�/�~�N�n����Mb�ɨ���#Aon�"�ږк30*�˽e����3�G�5M%�I,xr84�4��{�k�4)�<W
��)�����H5�&������:q	O߇���Ik������Ꮛ� �4�����?�{�?媁���l�v���c��� �G<^�36,�]���Ir|��'�+�ϓҾ����P�Z[=Q��v'�T�Ĵי��e�����v�񴲾	ڪ2N'�ھ5�&�/���CS�x{��P���)?*d�
0�+�ߎ�ܺ?���x{��ȎT���t�B�z1���U��'���^[CS[H��=*�=G�@�V!A#��i��UY��U��Ƅzk���|��K+�;ǭ�������|�x~io�,��X--�ES�]�(���Չ�� 
�N�$���Q�i��]*8dmSJi!h�Ta$q�
��夗�NJ�o�MQO����k-G�Qxr�8�o���	t��WE�H̋�`J�9�EzzT�l�x��Դn�_���W��A�����C���6�iZM����m�.�$�J�����b]��#�1#�׫[�}�o������#U��V���� �YB�)e�#�I�jFRV���)F�����<Ht?'H���[Y�ߺ��-��ne��8�ȓΑd�Ĉ|�R6�v!NO��Q�,M�h����,������+&��=�B ��N]��0�� 1_R����M*H�?��&��=9��0l��	���츧�x;@���.�t=6���J-���4x|�/.�+��f��$���F����i� �΅�Pצ�o�  �?�/���i��J������h��p��'�0v�q���![+2�_I���+}S��:�Z~�6���X��I�k[;�e4���s<2nr��2dm�ޱ�����N���'G���^u��P>ó+�Pp|��� a}Y�$��ɣ��m.��ص�&�ٙ�N>WfwbÒX�y4�:�W�����G*�y�,4� �� ��Vh�mm�+��F��&�t�/��i,��|�e�-��pa�!�~c�ܣ(����W�G��J�c�ҵ�� ���Q�L�1M'���Gp��1�s#0m�������S�Z:|��+a���m��� Z2p� xd�X�$𿁬�}*G�:M�׈n��D�L����y��J��V=r�	��U�1Jxw������?<E���{Q�-4�6[��E�wH��E�K�!�8�J�	/�ze�,v����޷�{�����n�L�+��v�����w��5��E�>���oB�������^��H�ՠ��VV�� ��?ϦB�Gf��2�dy^am���r~`H���_�~!��`6Z��r�v-ΘDw`�M�E9�,0]�� ��`~�E�+�Mt�� [���)sRv��^�hT��%'�<{�-/�wq@/t�+���+����������#� R�!�*g��M�Y�x�����\[�z�������i죹��Le��
���	1]%�ğ�W>�&��i��[�����P�>���
y��3I)����`#.�7�?��j:���H�O�o�x�3,��ku%�I�E��%�SH��D��nl�ii��5^_�������Q�Y�\��f��t��T��m���y��S3� 1)��d�Tt��Hԥ�s�x�����Z�O��P�e1�ڔV�0Y)0Q�к)�BW��}Ϗ������� O�T�B���]J�H2�Ȑ�m�d������Hbb(X����������e���<�4�4�"8Z��n�M�Y)��<�Y�-h�ܟ��ֆN)A^��z�v�������'���5{�m�����B���Ԥ�_,ϝ�����g1�z���K�xG\����v�$�%��n'�";.a�b�_242/*��m�}��AlMn���5�[\h:7�5K;aci��[Y�$�-�?��,Kt��l�6�l|ݝ��~\G�[G�F�6������+mI�DrH� X'f�6��f��Cr�����g
[�o=<�v9�������KOᩦO�e���;i��V�	��Ȯ�4G�fȔ��Bn�o�R�|ou��SK�縷��t�����ͷ[��1��!��=ˮ�$���W?-l|=�W�>!�O��[M�ִ�z��B�u;9��2�
�Cܯ�e�.~m�=�׀|1{�b�ÚMƮdIM��14��aF�
���Q`�-1�F4��(�� _Ռ���MN�_�� �y���+�?��xh�^]__^�铛�����+г��p�s"�Q�_��Mr?i�{���{� ���Zl�Z�N���R��f&1�\D�������=Mf]�m=�hdy��6�gGx�'u��4qƄ����x U[��ҋ�/ie�ϸ��D�����y��!O��S�[����� �B�C�'t���O��?�ӗ^#�.�o��W��-��׺��j�<V2,M���g��P�b� �f����g�މ��wG:]�զ�Dws��u,���lI
��k� IpZ8�J�9} � �)%��?�4f�x~��>"�ؗa]�+���q��?�q�|p�Фxc����I�%.eE�xW2HX	v�rj:���j�'����8�㴺��4o\iZr�}s=��i��ݛK���VGe��9 �%ĊZ%����s�w��i������{+�uT����(�U+ ��1�1	��� ���w9*�rk٫7ğ	���E�U���h:����(������k$%gR<ؼ��y��\�w��9�����H��T�|g����K	�_k�=��l��0���V��O6i"���y$|9�q��o�t��_�r>#i�md��	�ퟜֲA��KpQd��c�'��dB&�
�U#�Z^��Ί-ԋ���7���t�|�ymg�hdxf�����VV �:{��>�+�톭n6Gs�'cr@��s���v�ڥ����W�w1��\@��e]Xp�A�������n�SL�{%��,n�H ? �(O�s���T��*����O%���t������� �)���捧yX�=��y�����q�q�+�y���ʿ/�].�Fk��?l�r����ۛ�!X.���$.��&e�E�~o��8�,�5T�Gt�aH՘���#`z�8�'־.���)���k�z���6�J�tf�k[+��.��w�K���6�˱f���W�kN԰�]�穅k��Tkt� -������#���>#���w�t-"[��S�L�� !�2�8rHV��Q� H�������K���������5�x$q"�**�@  8 W��N�񆍡x�U�4�G]��]7��D/%�2J-e��[wI 3�����+��m�}�8q5�e}:7}|��(���(�� (�� +����� ��M�u��K�<��C'�$D�":�,�C)�� �E&�VeFN.�������7SL��6�'���+S&��	��܄���bH�SP��m�ï�����]�Q+��Q[y�)��!�|a�G�˸>�z����{���l�ͣ<���{�����rjzܖ���#�ĉ%ڐ�� �:.͢M�9 �b�U|�݁�~�>��ʻ�<@���&��Kl�Cj�o����G�6�\c�r����N�6���&�wR<�M��i�m��z���Om��[4��[O��y&��?�f�q�o��ݟ�2�:��� �~#�5�:k��OV�i�.���y��Y|�o5bY $(��l�۸�>�E5J	�m�u�4�{�yF��3�/UЮ�� ��B��%��Td���Kr�2���a��i ��U��Η�x�Mֵo��Z�������淑|�'Yc*�Hg`V�oRwe�j�Z(�4��W�<��w�����Ŷ�����;�&�j/���mgH��i�v�b3(v��*(��#h�:�%U�M݅QTfQE QE Aam�X�Y^��ygsC=��9Q�O�<k�� �z{~�s]���w~�o�5��?�ί��f��$H����b�'�@!�Ͽk�ϡ��������W����-D�io}�ӛi�x�!$m'�$��WR
9Ue8Շ2���S�V���_�� #'��t�t��M�[���ŕ��3붟d��+jH!p����)v��\&��� �`��W���im�n��&zs���{W�?~��#ď}7�~٥���GҴ�k%�[{5���'�{��ąb�خ����}�����x�������1�8Vv �GpMe8�Дd��7�8�	��]�#����!� �����j���u��|W�]�k�|9��s�k�[k��R�QD[�8tk�1�s�������j:������K�/v�ض3��g�+���P�6��\�� 	|�m� ������1��ͺi����f��d����H%V���TjҒ���:)ԭ)A� [�g���k��I� #�u����� ��)|��}��w���(������v�QE�QE QE QE QE v����� Q,����9'�����~
O`~����w���q[i6�Kk��S9`s��ݞx�;` (�w���� i6�Y��W��[��J���-�wg�z` �J�<V*u��v�?@�`)��I^Ovcj��uǞK���i�d��摍�� r01_>|R�C?�����-��V�L n�| 6�Ѱ98<�ӕSUҭ5�:{���u�$OЏ�A�rVx|T�I;�v5�`ib�խ.�������x%��Hf��6(�ȥYXA�A�Q���Q@Q@Q@Q@xw�K��<q�xo��/��/�����+=n��;N=B	c��K��Xѡ�� �`H�dR�+{�e\�n���Zv��(������YI�r���x��F3�8�Q��>fx���������<#�?x�S�6���Z�T��C�L�b-�M�ʫmBB�	$��(��qp����¬�Is+��� E���5�[� �_�XMk��N(d�{k��<�e#̅xd ��^#�^xf�T���Z���l�����'F�������m��c/��yx!���>�����!� �����j��{ᗈ&��t�x���R����a�2�4�n~�re/1�F㑣i\� F����%����鄡	�Kd��=��E}nڅ����c}���Dh���M�S ��_$�%�ݠ^�:�e�N���~ͧi���[C��ˊ5
���'
 �$����W����
(����(��(��(��(�������-�I��i�#yeL`ɴo��!��A�_1�!��� =�i��E��{��^ �rˀx��!��ҵ[MsN���t���w�*t#�r<�5���<�M�h�?E��!�������[��+X$�icR�$�U@�$���O<V�I4�$0ƥ�I*���I= ��ό �=�h�#y�c�k��B�b`�eT	$H��|<���Y�/O	M�O^���W���w��/�\�H���s1�8Oj��+�Ҷ��ٶ��QE(�� (�� (�� +����K�|:�V�d�Ky�iWW�$���⅝C A+���tu����Z�<�t_����(��������eu�v䌪Ƞ��I53�+��;s.m���<� G����z&�u�CB�ޗA���M��������r k�Wi�#����ګ�~|�º͖�����V���-`���
&���aV3	���D �6�N��)$��k�K���k����$���a��}-5�a����m���B�M�mB��c�,I��5�y�W��R�kP��ku�x��{#H���G��#3ʆ<]�&F%Nq���'�����@�y3�A;�#�$��.>��b���K���������6�{��$q"���@�x W=*� �+i���
8���o�}���9φ:�Z��-|]�x�����Z��kҨ��GT}���ld�(꫆�>5�C�w��wsk=�ZC�2�t�e���@ۤ�v*������Z;�}H�I�+_ ��*̂�(��(��+��~.��-�)5� 
ZCo�jV�9]W7��]����TI`�b�2����6��L����)ʧ�z��w�6�o�-CA:�� �zmΩ�\Asg?� �X��DS�ۆ��K	F?vw�N�����6������gf�2�wV����v���gM��9��)�w #/oO���k)�$�k<sC#�4l$����9Ѓ޼�ſ�H���A�R�V�e�M�Ϝ��K\����7.̏j�Dh���m�ؾ4�Q�N����R������0�N`�����B�m� ��H$
�k��=�T*��������N��o.%��|o�w.큁�y< ?
��c�?�/�<���j�}���;�G�H�r�g4qL��8,���U��j,����~8�,|K6���)��eg��y��jRd�#�R�HL�Ѩ�2�u
�6Oaʅ]%%������Z���@�>��M�j7���G��R�Ǚuoj�Qq�?�]���G����5&���Úߏ �����V�����&&�<��(Z����/�۾=絅�q{
�涇��^eᏏ�7��
��J�t�|Mj.��w=�fCλ���Pc���y �'�q�f�'NTݤ��(�3
(��
(��
�� �_��L�Zrj:~�yye{�hj����of���7I'�l��՗�Y_'����a.���6V�e���Hc�2-�H��7�������|� 7��[�5�y�]��W��+Z�M�G�Ɗ-��m�y���"0�-Ԣ9D£!�8U���V����u��	>i��7���N�e�� ��:�t�>�]�Ҵ�Ny4�[�&����Klh���p�@�6�`���׌t(f�&�K��C+)�A��������h����E�������}%����%��D���˹�$��}�M���5�Ѳ��Y�NJ���8��D��Aɻ�i*���*ڥ�}_�z���hxoUb�,.RFw>��
��vd$p>_a_|`�ό�kzM�r�K4h�c��k�II,̡��Y��I ����i�k:U�3:�u�����$dpk�-[M�F�ot��kY�h�*YX�# q�^v]5:R�� ��c9��W�"=4y7�5k� �_�Cm�P�S�,�K>!��L���*�#��'̱$���1��������u�湬�(�;��I�6���,����6ef��ۭ��)��D`�XI�E��ܼ�E{��k� 	���3~�jc�#Uo�	9o���;��N�����_?��+AF
�j��y�T��r�(���(�� (������Ƨ�/��z.�swc��j:\q_X��5��L-�\(R��	`!9ș7���]8��E�]��Xw	�n� �<�-� o�m�k�޸�.���&O��߲��)��9l��e�|H�w�|K�K?ĭ�j����i�Y�Ѱ�N��;)W���n�R�gLC i`o-k�5k��������j��Ƨ��u��ucj��Ʒ�a:%nk{E3�l'9��Ϋ)h��ǆ�5SZ��Ζ��m�ygy�Z�,vcN\�wl�ey�AS.����~\m����~
�<D5+[;����:1�7������vr��1�a]���q����O�5[�Vo�kqhQG�$��h�Vs�Xߙ���i$m�`���`�!8L����]ba��C\��5����]�Ki�ᕎ����L� A"H�p*�e $�J\�?�Rx�E�S{�� 3���.���h���E"Ѯ��t�3$����ŉ��g�%�d�c�`�9��b��v�+�Lݯ�\�w��%%��+if�0����$�󍯄�"�;��m��}��^#�t�:�V�廋T���**#����� k��=�Q񦹫�n��� �;q�x�P���#� D�y�1�f�����9i�D�~TQ�+8u�����=>��w7�|}��N��U�Y����Q�����I ��Po��Ϝ�}ڞ'�w�� ��u�Y=��'�|��aY�ݻʙQ�My� e��ɯ��Ŀ�~�/�u�oD�������t�;�/����(��Sm(�'���E�F�Y�����#����?�� ���<ikh���u[f�aj��������ڰ��0�:m��䉕*я;���� ��O��Mf]TiR}�K��,on
,�u�2��j�{xd!@���0:�W��C�?��-e��&vv��`����w�~�?{<̻��dm�A���m�]�e֮m�4+��Z�AWK1��&pv���!l`e�ۘ�<9��K��J���ĺN���+&�>�^$&�Pi#gk�ڲ[ق�$�l-ā�l��R�&�.Tf�̪]Z�W��G��	|��sD���]>��9P�kI�۠X�M� �WRpX�d���W�Z��|+�x�i�������巻��#�پ�[1u��M�# �}'��/���~��^���a��\���]��e�/�YJ���Y]V��mR�F�b����	�J�M[�{��
�/�u����� ��i�4�ZxzT����9����<0�-��7�Ғ�c����SWG%Jn�I�QVdQE �$�!��ⶩ�x�S�ޕ��~��J�ݩT(��[�ڈ �z��pN`��u�:��_ؓk�~��j�/�bԢ�kk�,�Gr���ѣ��yȑ���+�����k�Ϩ���͌w����J��-5�2���Gpش�pwyȤ����fz朔���o�~����(Cک8����oӷ��X[iv6�VV�Y��F��o�$Q�EQ¨   
�� ٯF�c��α7�"Z������g)�C�^z
�z���� �Gn�_̒�?�09ؖ|�sq�c5ǘ��Ⱥ����Qu1��?����_:�о�N�$Z�a��PP�1�ʊ0P$�~¾��Ǟ��~�� ��}�����9S��H�Xw�	[�UR{lϨ�᾵A�o��??>4xoN�<+%δ�%��lc���?�'���C��%u��]'2eW+��������MkW>���n�����4�T�mד�1�q��H�hÖ(�=fx%��Hf��6(�ȥYXA�A�_|M𮽨��M;�6]�t� �Mo�b4c~��O���K����f ��Aկ��hITJ� �W���:ub�7o��[���>���_�:��|!i6�o��տ�#�kz�M�4`#]�mšI3*8F�@�=UuE�+��Qqn,(��K�~���⾎��Ԯ�k����c�{�e�yu1x����������|��N���NǶ�_/�gK�+��u�aҥ��� J1��4��>z��k$����k�����2��ď|R3�[����Fa�^�~o�l�1s�HZ�5�@�c[��!U�1������� ������\�����CQ^�� �ڟ��B.�Q� ��z�L��9'���r9{heYv��Ŏ/1��B�-k|,��7�;�Xx�X�RCg=��/��F�-Ǜ�o�|�r���:�*�d�ʖ� �r�nJ��Ǵ�_2�z��W���"t�{�����"�/o�ή�r�"�z��,�k��$_2m��I����]���6V�����T�S��tg""Z�%�I������̱�_#%]=�*XV����_��r��U�w��'��=� ���� ��+k�cѐ%�ek�mfw2F3/��+#�� �w��CĿ5/|?MN٭4���]��{9��C)�X��ž�a�d?���R��'��/�-/���xOC���{���~�y���X�^Z��Z�T��C��ʏAZ��^	׼{�o���Z��mu+?K���D��kq䮯H��UZ�K?J8
k�l����[�/�]�3[�m�8��L��R��{o��g�J�FR�_1v���Y��R�ԥ����֍���=l}gE|�.���Z�s�i"�C5������뢤ήb,�Z�R|�#�� n+���K�VV����:F�y�/P��إ��m*[�A�;ܪ@\��,�T�8O��c�����Ϭ诖|7�?��f����|yxST�[S5Ɯ��a���&)C0R��D��2����/>@_�=Z{z)$�t�%�1�ɧ�l�5x����ŖX�۸)k����I�̷���6��g�n�s��!׎�j'�G�h���ؑ��&gT7A� (M�J�y���{�Pj���a�Yxb_]F�������5������%uk��r�^5���b={e����g��O����_Ǘ��߄V����o���jz�2Aa�G�+X]b�Cȱ�|��d���$m�L���|Tҟ����|/�K�&���c�����a�(����I�����EG����>��ȍ�h���e�o�_�=K�ZTv��[E��~��{+I�»��^K���o���um�,wyTPi>�,)J�\���������x��Z�����CJ�����6�������Q����Kig�H��Ơ���T�9+�����x�œh���+�~�q����_.-�'h��|ˆ+��R\���;B���ݍ���&��ڌ_j������4R	���m/��h���ET"��Lc��pR������GMj�0�+O����_'c��/�I|K�kI�u��Yn�r>e9�s�2X2��<W���|�o�"�ϋ��oqqs�pˑ�FrW�9����o[�Uv�h}�Y���_w�
(��X�?����q�]>$Ky�%�Q��BN%8���6:�5�w�� �c����Z>��ܮ��=��5a�p�C����1d+"�����Zk�t��%ͤ�H��Ѓ����~&x_ k��d{�	��m;)�pQ�0Yx�;<g��8�V�{�����pr�S�4��_�g�:u���C�T���3��F����B�D������>�f�7S:�2I$��$-��K���V�<�K��>�C��ڭ�]��e�U$��fy_�y0����[/���~ҼK�|<�o�]�u�\Ũ�i��ƫk	/-�SD��� ��H��9�?�îx<)>������}�v��h�h��-��]Y�S<���y��k�3J�u��%�]����������o}��UQ]�ex�z���-F��h��͕4�T�d�0@2}�j�E	%�m����(QE QE QE QE QE QE QEQ���/isj��E�[A!ٙ�*""����UQAffUPI��cI�dr�m<A7��J����vzޕ�U����������n��))@�F�� d�do Ѵ����h.~�w.�?�t�Yŧj����u	$�1%�嘻���غ���<�^�������|S�Aw&��=F�M���M�M�H�=�̳����$�dǕ#\�,��O��_�9�j�日Eg��4�R�6�w��:!;ci<�̅�h_qPG��ji� _��zjUN���]t���kS��J�%��|Y���}I��0��J�!�B���CW#�	����V�U�y^fZY�X�rX���$��������!�æ��P',����ݏv8�@` +v'�C�����:���T��^��Y�EW�tQE ����x�@��.��I�V]�0v�9�}FFA��٢�2qjQ�(�qq��g�>'�ơ�bm7R�ʝ9V^RE��{���\���]'F�u�^��(5=fH���2\�X�O�(F %�2�O��~��GHĿg�mw5��N̜eXt�s�`�A�����<!�M��P�S�*��H��Ou8�`��+�0���"��/���� ��o��}Fy��&���O��~���$���f�s{~t�qpȲEi��K3F���D����������ޭk�y��}Q��I��0�)�HѢ@Ī�Ip��
P�7㟂�x�Y���F���cW����i��q(�G����P��pfo�������h!�[�rGs�[[۹�cҬ34wV/��.�e�d�"{h� �"���N��Q)l�?��� �-�4iԤ�ջ�=:i����������������R��u{o�Y��<K=���,q��襾b�,0�Ǡ5��e��y�-%.�ES$(�� (�� (�� (�� (�� (�6_�>����<E�j^.1��G���3C��H����AR�W![cc�u� ���� ����hVq�Z֯m��Rx~�w�Yda'�-X,���/�U'��XG��=I}�o����zw��!Yi_<K��ԃE��%hr����VX����.��Gϑx�G�t�.��x?U����S�n�����V�#y	i>��u���wp���*v��o������L���!��_Y���x�Hb>ũ�,�JyBG�#��M,� �|�od�>xw�ڤ7�V�a�}��}F�{[<�_�{y$h��3"�h�Q�
H8k]y_ד�Οw���v�~��"���7���ݦ����;3W����zTzh7S�ח&������A���KJҮ��F��v�Iԟ� �$� $ѥiWz���sw;l�$�O� d�x k�O�?
W�)=���s�Φ&hX�Qǐv�@�$I��εh�"�wodo��O0�RV�ѿ�����o�X<���1���=��jx��d�A����5��E|��*�r����t�J
VH(���@��( ��( �/x/I��j��o���26�"$c*#��H�ETd����Ȝ#R.3WL��_�o����i�!����ddg*��}���+�WJ��4��/�K�I�d�?B?�� ^㯀�<f���K�����/���0$���@ɯ����Qr�����vS:M΂�{u_�|��OiZ��]o�h��[[XxgJ%��nu)a��yK/�	.+�d� �C{��F����O�R]KU��#�{�&T�Ңy2��aP�H���`}Xz� �?�t�贻��=F���}m��є3*eFXc��p-(x#��|��� _՗��F�y%+� ��߫0��sL���di�j�-֩�k�[�p/�M��|�D�E�h����wP�����O	|1��� ��]���.E���X����8j.F���s��|���_���D��Yt���3][ؓ��q,��y�9��q�Q�F�ry�~/x��n�{��gO�oh)�%����-���o��S�G���,W�
���q ��PW�� ^A��J��¼� �>�.���h����m.KG�m5]:}�U��42a���RA�PE^��>|C��s��|{��$����Ի�Hӯ���fH̕�g%(>�(��c"v���$�U״������ư^��������ǔ���K��/��wS�$J�E���Y�p�����O%S�;7o���K��Ey���OI�#@�/�uO�Q�֥<�^��a���[�m��d� �YT�̜+f�/�N�5� 	?�#��_��#�}��y��wo��7O��J�N/��*S������Es����o_=��������gX�W2�S4x� Ys�șP��N�e<7���0�_L�5��IVC��G#��0�Ja��/�$�3�ƎX*�#
�9㦻���_u�vTW�|T���k��O�|Wc�j%X�_�ZK5������&��<�G�[rIu��*��Y��E��zd��K��,�E�{{Y��1�y^�~��a�$��O]��=�u���MVz_K��=:�� �ǂ/� |.ִ�)�:��Ϸ�K�`���-i)�X�ɾ&�&��5��~|.���Mm5��e�xFMz�� 
��km*�%�Ȓ*��6�fǹ|-}M�	�.�ai���6�6Me�I]m�mݙ�� ��Lw!b���^6ѣGNXf�y=��� �|���˻��>���{��GN�� u��kp���5��W�y�5���9P7��O�i�X[x�ƺͿ�>j1x{�~9Җ�S���&�}>�(��g�ݦT2ʍ���V�_t��?����.�Eo���_��������k:i�x���	��Q����n9'�������i���1Q�,�߳��vz���exO�v�𮍠Y<���VP���dd�)b ��8 g����~ռk|��U����2��8�8���d��u��	j^,H��&}/IuY#|,�O���� ��;�����1�?�<:n��r�ܼ����c�� ��8�Q\���;�y]LK�����ٕ�_��O��G�#��G=��~Nrp3�\���H�utQ_59ʤ���ϵ�N��d��(�4
(��
(��
(��
(��
(��9O�1�� �7I}i�^�}�"9�������b�;�� �A���X��ݘ�;T"a�G1rz��Kp	8��(��ʴ4N�<�N]C����Z�O���Ѽ3F�9�+�==�:�7�>�|Wj-�k�c_�\aӐN�e�ќ�s^k����]��f��\i����M�@'��� r9,O���*R�տ�����I�/�� ��|yu�NҡХ�{E�k�
K���c�[ �N^�m�X��ϵ�(G�2�U(p��W�g����^������!�M+���v��2ʖ��5(?z�$���N����ŶW����9�-�]��_3g\��Cӊ�'�}�{i��?�������8`#�댰��-}������������ϛ�!�յm_�2��� �Q���A7��6��O�EnR��݂�	X	.���*FQPW����O���&zW���V��ŵ��A�SL��I��zH��2��7;�}��R�w��� ���q����>x�[���z'�~�kpkw�7�4��^mN��;��1A�QZ�,�S��kP���*��7��x����6m4�ό��/&�S.t���_-nw��P7F�V�4T�����H�b�'{/ӯ���5���%�SU��x�Ѿk:�����R���-�w�Gqу��@�.�Y6|��z��A��{�~��cci�[��$Q�������I+��ϙ���a�+rȬ=J����B��E�Gg#+)9w��M�����9�-���Ksp�I���{�y�Lq֡���_6i���B/䭿���y������R�o�H&�x�+L��y�".O8U ���4oٮ�6����.c���G����nQ����+Ӽ7�}�;Γ��i#�t�/!]�Km�A�q��W-Lƌ>��M���Q�� _3�_
|�'�gkG�����!F�3�3�1���n���=�� yS��Z�a��tma���� ��$n5��^5lmZ�^���<6Y��kk��(���=`��( ��( ��(������ JFIF      �� C 


�� C		��   " ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��(������ JFIF      �� C 


�� C		��   " ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��(������ JFIF      �� C 


�� C		��   " ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��(������ JFIF      �� C 


�� C		��  � " ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��(������ JFIF      �� C 


�� C		��  � " ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��( ��(������ JFIF      �� C 


�� C		��  V K" ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? �S�����������:���:��������/x�➗��Z�J��Rյ{��ج4�>s��c#���g��2�|o����;,�'�d�A������|�/�	%���œ��Z=�?`���M�5�b��ۺ� v��U���^-���mv?����}\��2EP���"gʛzn���T���ri${�1��|{�cK�ͦxw��|ckiv��z���*��S��|����S��� ����!.��D���c{a��Z�2Y���$�K�"�����i���I^�;����4�Y����ij�v7<G��C����Y�������ai�Z[JX�&Fo\� ��VW�jV�\[ʓ�*����WSЃ_7|iԴυ_t� �R��²�Kl�_3-'^���|�W�K�����t�lt]WI��J��;[{�g��0���՗���pM�PC2\ƒ���eެ���9���J�U�˨LMĻ��c�st�$Q�v����_x�ŷ�;�M�~�n��ˉ�o&=�,C�J����k��-�Q$�� ��d��� ����}k��>
C�����^�h4_Z����_�;�D��$�����2v4�Nud�v� M��>��-��I��zo�,����-CT����Ka>GmꍶO�m7���M�S�������t�/	y�[��|����+��ƿ¿-c�w�z�����ZD��iaw�	A�d�N���MZB����q%Ǜ�&�yo-��~��3�+C�M��&�]:����k=;T֣��E�P��ߕ��+򍣌��� ���SFQ�����٤�I���_���ÿ���mL�_�4�����F���Sd��۳�8��i2��$���y�xo�>x��?m��
|.���k;Wk��1oᑉ�|�o<ya���x�H�e�� ZѼ7�j}\��b���{_\ϳ������n;|���V�n��h����*ҥ������FV���S��P�FJ�[Ϩ��M��ZS�75/�&�^��}���/�Z}���|S�Ƈk�"-�K���c�47��)]��ޡ?�nڙ�^�h����P�c�C�2��,SB��Ȏ����5��j?�!h���4ۨ��$Z�&�'�ŝ�r]�%�����7�+E)T�>�M�k���
'��	[���O^������	b���41��X��/�H߼�iM�}�:�Y��q���j?Z���{%m��e���\�� ����zv���ג��)�V�����;�~�ww������x7�O����o\���=��u�6���q�u�evVV��.����������ߵ��.���*���to
k֗v"�d[�{�L��Nc�$1���oz�+�y'�A�m�<cw�8�	t9썅��R��*�,-�F�x2�ɥ+[S�9�g�v��{�b���v�
 ���<w3j��ޒ��v��Hm�bD���QF�B{⼇����5�?�t������O�Γo1��������_�z~����Ŗ�0^X}m �V;�1�k����_#��l�|}2�\�$��ɩHש���@ɷ��w����5c
�'V�u�_�o��<w�O\j:i:u��	c�k���k�ʣ=Q���Y����_x�࿍O����{_�Kw��sFp�[ië}��g�hm{��&��-pI�[U�� �Iu�O?�k����B̸U��v�^v��k���_����t�4�S�R��v�n�b��T�d����V�ˉ�<����G� ��k(�2mu[��++���L��?��]t�[�#����Ǟ����0����� <�p��u�������<;��������hz�Q�6q������� �̮�������<� �f��~Ȟ'e��|8�FE��DUژ�$���b��Ğ9��3�]^]/��е��Hw@b��������G��e7[��2��ץ)F��f�J�+��Σ
��))j�(`��C�����?
�����S�5�ٮ/�kˈ��}�U�!��y�e��)�������q_�Y���J�U����o��#g�:m������WU�%�����?���������� �緓�r�s�����W�7D�~�^��'~�S�k�&��v�$:to$�pM��䴘��w?v�^{���s��,�X��x�{�>ק^-������FY���u�G��i���>0�ռ;�yt���[���ⶹO+�P��^Bg�~_��/��Y_|C�����i��Ai}-�Z4�m	1T�#Ʋ�R�W~ߕd�Kㅯ�r�K�y��Gu$���[7��(�Ѽ/�^Y��h=kǖ�����S�FGi��������x���M{�	>�/��o�ͦ����g=��؄6�l���M�.�[> ����۳Y��$� 
5MǇ�ЯlZ�Oݏ�	L����}ݝ��5�xG���߄ �V�ᯱ����������-�ZOp���"l�~g]����Y(�d�e����ؼM:TjԦ�*�MN.ܰ������v3?f�F{?��M�Sl����?��|�I\'�����Ǿ2����˛��'Ŗ��w�«٬�n$,��[_��­�|��|�YM�&=��>���N�k�D�W�H���b�j��h�^x$�5�����\����"o+v� G��,c��8m�Z������d�pS��uk||�my���h�F�Xcp0T�y7���x��ׇ�O��o�$Yc���ѭ%�L��6
�EV�k��ڵ��h����
��&��Zj�O�0�U}{��R��4��u;{y%��,f�P��{��]���zf�9�m�G�:��u׼/��Z�~��5��Ko� (�N��T�� gVܪ�{g����گ᷌~-�,>�Uޝ��7��\]j�	�(_�V��V"O68��;���w�2�p��?b�oD�=�Ӥ��^2��e��P}��f��� c�� w*�m4����#鲅B4%�%N�i;��՚�&�b����u�!���qk���k���s�kV���i��gm�d�Kqq���?�6�?�G��I|Eo����R�G��m;e�%?8�)�\'�?fϏ�9��j�τ-�񝕅���j7����H�<��#e��/�����7��w�4�'ŒA�j�������1m����wvZ!{�_��o�j(U��v��V����m/$|w��p���llu�㴃�U�gؿ�H��:|O�W�����ZTfc$��F>c�|�����v>"���I���Q�_�N�-6&i>I$V�o��ߖ���'�=W�`��'���>_�ݙB�����Z�|���o�~-h����3���%��{j�c_&�=��H�W�#V��2oy�������ǩ���x�x��� Ey��F}66��C�,[ك���O�;ڻ_��.x������z.���xZ�Ñ��R���1w�L~\�:���HG������]+P��>#���h���[k덂]�y�V��9L���ڳj��X9P���n�v���}���m;���^��D��&��i���b���I{�cX��
ɍ\E�6�֖J��{_|%��>/�ǟ5WĚm���]&�K����4�4�6t 2*}�l�u��}��z�^ڣ��)ҍd�J-5�om4�դ��EU�HQE���wO�������s�;.ɓv����'��k�E QE QE ��    ��E ��E  |�� ��� ``` ����                   Texto circular���B���B���E���E      �A��� ��� ���         ��� ��� ���   @        B   @]   Aplicaci�n de Manejo y Consulta de las Referencias Bibliogr�ficas de la Traducci�n del SWEBOK         Arial  �A             Texto  E @�E �E  �C     �A��� ��� ���         ��� ��� ���   @        B   @   Trabajo Fin de Carrera         Arial   A              Texto #2 �E ��E �+E  �C    �A��� ��� ���         ��� ��� ���   @        B   @   Manuel Monge Mart�nez         Arial  @A              Texto #3 P�D ��E xE ��C     �A��� ��� ���         ��� ��� ���   @        B   @,   Ingenier�a T�cnica en Inform�tica de Gesti�n         Arial   A              Texto #4 ��D @E  �E  D     �A��� ��� ���         ��� ��� ���   @        B   @I   Escuela T�cnica Superior de Ingenier�a Inform�tica
Universidad de Alcal�         Arial   A              Imagen �2E �(D 0rD ��D        ��� ��� ���         ����                   B                        K   V       ��� ��� ``` ����                    �e�E�e�E  ��� ��� ``` ����                     ��� ��� ``` ����                    ��F��E  ��� ��� ``` ����                     ��� ��� ``` ����                    